package rd_dma_regs_pkg;

parameter RUN       = 0;
parameter BASE_ADDR = 1;
parameter SIZE      = 2;
parameter IRQ_EN    = 3;
parameter DONE      = 4;
endpackage
