package rd_dma_regs_pkg;

parameter RUN       = 0;
parameter BASE_ADDR = 1;
parameter SIZE      = 2;
parameter DONE      = 3;
endpackage
